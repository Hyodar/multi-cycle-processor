
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package unsigned_array is
    type unsigned_array_t is array(natural range <>) of unsigned;
end package unsigned_array;
